`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    08:12:57 10/19/2016 
// Design Name: 
// Module Name:    GenColor 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
/////////////////////////////////////////////////////////////////////////////////
module GenColor(
input wire col ;
input wire row ;   
output reg  
	);

if (row <= 200){ 

}else  if(row <= 400){

}else if (row <= 600) {

}else if(row <= 800) {}

endmodule
